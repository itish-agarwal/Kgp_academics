`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Create Date: 12.10.2020 14:35:47
// Module Name: 16-bit Arithmetic Logic Unit (test - bench)
// Project Name: Ass_5_Grp_6
// 
// Assignment 3 - COA Lab
// GROUP 6
// 18CS30005 - Aditya Singh
// 18CS30021 - Itish Agarwal
//////////////////////////////////////////////////////////////////////////////////


module ALU16bitTB();
  
  reg [15:0] A,B; 
  reg [3:0] S;
  reg M,cin;
  
  wire [15:0] F;
  wire cout, is_equal;
  
  
  ALU16bit myALU(
    .A(A), 
    .B(B), 
    .Select(S), 
    .Mode(M), 
    .cin(!cin),
    .F(F), 
    .cout(cout),
    .isEqual(is_equal)
  );
    
  
    
  initial
    begin
    
    
    $monitor("A=%d, B=%d,S = %d,M = %d, \t F=%d, cout=%d",A,B,S,M,F,cout );
    cin=0;
    
        A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0000;M = 0; 
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0001;M = 0;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0010;M = 0; 
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0011;M = 0;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0100;M = 0;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0101;M = 0;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0110;M = 0; 
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0111;M = 0;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1000;M = 0; 
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1001;M = 0;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1010;M = 0;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1011;M = 0; 
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1100;M = 0;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1101;M = 0;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1110;M = 0;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1111;M = 0;
    
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0000;M = 1;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0001;M = 1;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0010;M = 1; 
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0011;M = 1; 
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0100;M = 1; 
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0101;M = 1;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0110;M = 1; 
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b0111;M = 1;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1000;M = 1; 
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1001;M = 1; 
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1010;M = 1;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1011;M = 1; 
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1100;M = 1; 
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1101;M = 1;
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1110;M = 1; 
    #10 A=16'b0001101000101101; B=16'b0010011101110011;S = 4'b1111;M = 1;
    #10 $finish;
  end
    

endmodule
